//
// SCARV Project
// 
// University of Bristol
// 
// RISC-V Cryptographic Instruction Set Extension
// 
// Reference Implementation
// 
// 

`include "fml_pack_widths.vh"

//
// Checker for bit packed multiply instruction.
//
`VTX_CHECKER_MODULE_BEGIN(instr_pclmul_l)

// Pack width of the instruction
wire [2:0] pw = `VTX_INSTR_PACK_WIDTH;

// What we expect the result to be for a pclmul_l instruction.
reg [31:0] expected_result;

integer i;
integer j;

// Partial results
reg [63:0] pres [15:0];

localparam SHF = 0;

always @(*) begin : compute_expected_result
    
    expected_result = 0;

    for(j = 0; j < 16; j = j + 1) begin
        pres[j] = 0;
    end

    if         (pw == SCARV_COP_PW_1 ) begin
        
        pres[0] = `PW_CLMUL32(`CRS1[31: 0], `CRS2[31: 0],32);

        expected_result = pres[0][31:0];

    end else if(pw == SCARV_COP_PW_2 ) begin
        
        pres[1] = `PW_CLMUL32(`CRS1[31:16], `CRS2[31:16],16);
        pres[0] = `PW_CLMUL32(`CRS1[15: 0], `CRS2[15: 0],16);

        expected_result = {pres[1][15:0],pres[0][15: 0]};

    end else if(pw == SCARV_COP_PW_4 ) begin
        
        pres[3] = `PW_CLMUL32(`CRS1[31:24], `CRS2[31:24],8);
        pres[2] = `PW_CLMUL32(`CRS1[23:16], `CRS2[23:16],8);
        pres[1] = `PW_CLMUL32(`CRS1[15: 8], `CRS2[15: 8],8);
        pres[0] = `PW_CLMUL32(`CRS1[ 7: 0], `CRS2[ 7: 0],8);

        expected_result = 
            {pres[3][ 7: 0],pres[2][ 7: 0],pres[1][ 7: 0],pres[0][ 7: 0]};

    end else if(pw == SCARV_COP_PW_8 ) begin
        
        pres[7] = `PW_CLMUL32(`CRS1[31:28], `CRS2[31:28],4);
        pres[6] = `PW_CLMUL32(`CRS1[27:24], `CRS2[27:24],4);
        pres[5] = `PW_CLMUL32(`CRS1[23:20], `CRS2[23:20],4);
        pres[4] = `PW_CLMUL32(`CRS1[19:16], `CRS2[19:16],4);
        pres[3] = `PW_CLMUL32(`CRS1[15:12], `CRS2[15:12],4);
        pres[2] = `PW_CLMUL32(`CRS1[11: 8], `CRS2[11: 8],4);
        pres[1] = `PW_CLMUL32(`CRS1[ 7: 4], `CRS2[ 7: 4],4);
        pres[0] = `PW_CLMUL32(`CRS1[ 3: 0], `CRS2[ 3: 0],4);

        expected_result = 
            {pres[7][ 3: 0],pres[6][ 3: 0],pres[5][ 3: 0],pres[4][ 3: 0], 
             pres[3][ 3: 0],pres[2][ 3: 0],pres[1][ 3: 0],pres[0][ 3: 0]};

    end else if(pw == SCARV_COP_PW_16) begin
        
        pres[15] = `PW_CLMUL32(`CRS1[31:30], `CRS2[31:30],2);
        pres[14] = `PW_CLMUL32(`CRS1[29:28], `CRS2[29:28],2);
        pres[13] = `PW_CLMUL32(`CRS1[27:26], `CRS2[27:26],2);
        pres[12] = `PW_CLMUL32(`CRS1[25:24], `CRS2[25:24],2);
        pres[11] = `PW_CLMUL32(`CRS1[23:22], `CRS2[23:22],2);
        pres[10] = `PW_CLMUL32(`CRS1[21:20], `CRS2[21:20],2);
        pres[9 ] = `PW_CLMUL32(`CRS1[19:18], `CRS2[19:18],2);
        pres[8 ] = `PW_CLMUL32(`CRS1[17:16], `CRS2[17:16],2);
        pres[7 ] = `PW_CLMUL32(`CRS1[15:14], `CRS2[15:14],2);
        pres[6 ] = `PW_CLMUL32(`CRS1[13:12], `CRS2[13:12],2);
        pres[5 ] = `PW_CLMUL32(`CRS1[11:10], `CRS2[11:10],2);
        pres[4 ] = `PW_CLMUL32(`CRS1[ 9: 8], `CRS2[ 9: 8],2);
        pres[3 ] = `PW_CLMUL32(`CRS1[ 7: 6], `CRS2[ 7: 6],2);
        pres[2 ] = `PW_CLMUL32(`CRS1[ 5: 4], `CRS2[ 5: 4],2);
        pres[1 ] = `PW_CLMUL32(`CRS1[ 3: 2], `CRS2[ 3: 2],2);
        pres[0 ] = `PW_CLMUL32(`CRS1[ 1: 0], `CRS2[ 1: 0],2);

        expected_result = 
            {pres[15][ 1: 0],pres[14][ 1: 0],pres[13][ 1: 0],pres[12][ 1: 0], 
             pres[11][ 1: 0],pres[10][ 1: 0],pres[9 ][ 1: 0],pres[8 ][ 1: 0],
             pres[7 ][ 1: 0],pres[6 ][ 1: 0],pres[5 ][ 1: 0],pres[4 ][ 1: 0], 
             pres[3 ][ 1: 0],pres[2 ][ 1: 0],pres[1 ][ 1: 0],pres[0 ][ 1: 0]};

    end

end

//
// pclmul_l
//
`VTX_CHECK_INSTR_BEGIN(pclmul_l) 

    // Correct pack width encoding value or instruction gives in bad
    // opcode result.
    `VTX_ASSERT_PACK_WIDTH_CORRECT

    // Result comes from the PACK_WIDTH_ARITH_OPERATION_RESULT macro.
    if(vtx_instr_result == SCARV_COP_INSN_SUCCESS) begin
        `VTX_ASSERT_CRD_VALUE_IS(expected_result)
        `VTX_COVER(pw == SCARV_COP_PW_1 );
        `VTX_COVER(pw == SCARV_COP_PW_2 );
        `VTX_COVER(pw == SCARV_COP_PW_4 );
        `VTX_COVER(pw == SCARV_COP_PW_8 );
        `VTX_COVER(pw == SCARV_COP_PW_16);
    end

    // Never causes writeback to GPRS
    `VTX_ASSERT_WEN_IS_CLEAR

`VTX_CHECK_INSTR_END(pclmul_l)

`VTX_CHECKER_MODULE_END
