//
// SCARV Project
// 
// University of Bristol
// 
// RISC-V Cryptographic Instruction Set Extension
// 
// Reference Implementation
// 
// 

//
// AES SBOX function
//
function [7:0] sbox_fwd;
    input [7:0] in;

    case(in)
        0  : sbox_fwd = 8'h63; 128: sbox_fwd = 8'hcd;
        1  : sbox_fwd = 8'h7c; 129: sbox_fwd = 8'h0c;
        2  : sbox_fwd = 8'h77; 130: sbox_fwd = 8'h13;
        3  : sbox_fwd = 8'h7b; 131: sbox_fwd = 8'hec;
        4  : sbox_fwd = 8'hf2; 132: sbox_fwd = 8'h5f;
        5  : sbox_fwd = 8'h6b; 133: sbox_fwd = 8'h97;
        6  : sbox_fwd = 8'h6f; 134: sbox_fwd = 8'h44;
        7  : sbox_fwd = 8'hc5; 135: sbox_fwd = 8'h17;
        8  : sbox_fwd = 8'h30; 136: sbox_fwd = 8'hc4;
        9  : sbox_fwd = 8'h01; 137: sbox_fwd = 8'ha7;
        10 : sbox_fwd = 8'h67; 138: sbox_fwd = 8'h7e;
        11 : sbox_fwd = 8'h2b; 139: sbox_fwd = 8'h3d;
        12 : sbox_fwd = 8'hfe; 140: sbox_fwd = 8'h64;
        13 : sbox_fwd = 8'hd7; 141: sbox_fwd = 8'h5d;
        14 : sbox_fwd = 8'hab; 142: sbox_fwd = 8'h19;
        15 : sbox_fwd = 8'h76; 143: sbox_fwd = 8'h73;
        16 : sbox_fwd = 8'hca; 144: sbox_fwd = 8'h60;
        17 : sbox_fwd = 8'h82; 145: sbox_fwd = 8'h81;
        18 : sbox_fwd = 8'hc9; 146: sbox_fwd = 8'h4f;
        19 : sbox_fwd = 8'h7d; 147: sbox_fwd = 8'hdc;
        20 : sbox_fwd = 8'hfa; 148: sbox_fwd = 8'h22;
        21 : sbox_fwd = 8'h59; 149: sbox_fwd = 8'h2a;
        22 : sbox_fwd = 8'h47; 150: sbox_fwd = 8'h90;
        23 : sbox_fwd = 8'hf0; 151: sbox_fwd = 8'h88;
        24 : sbox_fwd = 8'had; 152: sbox_fwd = 8'h46;
        25 : sbox_fwd = 8'hd4; 153: sbox_fwd = 8'hee;
        26 : sbox_fwd = 8'ha2; 154: sbox_fwd = 8'hb8;
        27 : sbox_fwd = 8'haf; 155: sbox_fwd = 8'h14;
        28 : sbox_fwd = 8'h9c; 156: sbox_fwd = 8'hde;
        29 : sbox_fwd = 8'ha4; 157: sbox_fwd = 8'h5e;
        30 : sbox_fwd = 8'h72; 158: sbox_fwd = 8'h0b;
        31 : sbox_fwd = 8'hc0; 159: sbox_fwd = 8'hdb;
        32 : sbox_fwd = 8'hb7; 160: sbox_fwd = 8'he0;
        33 : sbox_fwd = 8'hfd; 161: sbox_fwd = 8'h32;
        34 : sbox_fwd = 8'h93; 162: sbox_fwd = 8'h3a;
        35 : sbox_fwd = 8'h26; 163: sbox_fwd = 8'h0a;
        36 : sbox_fwd = 8'h36; 164: sbox_fwd = 8'h49;
        37 : sbox_fwd = 8'h3f; 165: sbox_fwd = 8'h06;
        38 : sbox_fwd = 8'hf7; 166: sbox_fwd = 8'h24;
        39 : sbox_fwd = 8'hcc; 167: sbox_fwd = 8'h5c;
        40 : sbox_fwd = 8'h34; 168: sbox_fwd = 8'hc2;
        41 : sbox_fwd = 8'ha5; 169: sbox_fwd = 8'hd3;
        42 : sbox_fwd = 8'he5; 170: sbox_fwd = 8'hac;
        43 : sbox_fwd = 8'hf1; 171: sbox_fwd = 8'h62;
        44 : sbox_fwd = 8'h71; 172: sbox_fwd = 8'h91;
        45 : sbox_fwd = 8'hd8; 173: sbox_fwd = 8'h95;
        46 : sbox_fwd = 8'h31; 174: sbox_fwd = 8'he4;
        47 : sbox_fwd = 8'h15; 175: sbox_fwd = 8'h79;
        48 : sbox_fwd = 8'h04; 176: sbox_fwd = 8'he7;
        49 : sbox_fwd = 8'hc7; 177: sbox_fwd = 8'hc8;
        50 : sbox_fwd = 8'h23; 178: sbox_fwd = 8'h37;
        51 : sbox_fwd = 8'hc3; 179: sbox_fwd = 8'h6d;
        52 : sbox_fwd = 8'h18; 180: sbox_fwd = 8'h8d;
        53 : sbox_fwd = 8'h96; 181: sbox_fwd = 8'hd5;
        54 : sbox_fwd = 8'h05; 182: sbox_fwd = 8'h4e;
        55 : sbox_fwd = 8'h9a; 183: sbox_fwd = 8'ha9;
        56 : sbox_fwd = 8'h07; 184: sbox_fwd = 8'h6c;
        57 : sbox_fwd = 8'h12; 185: sbox_fwd = 8'h56;
        58 : sbox_fwd = 8'h80; 186: sbox_fwd = 8'hf4;
        59 : sbox_fwd = 8'he2; 187: sbox_fwd = 8'hea;
        60 : sbox_fwd = 8'heb; 188: sbox_fwd = 8'h65;
        61 : sbox_fwd = 8'h27; 189: sbox_fwd = 8'h7a;
        62 : sbox_fwd = 8'hb2; 190: sbox_fwd = 8'hae;
        63 : sbox_fwd = 8'h75; 191: sbox_fwd = 8'h08;
        64 : sbox_fwd = 8'h09; 192: sbox_fwd = 8'hba;
        65 : sbox_fwd = 8'h83; 193: sbox_fwd = 8'h78;
        66 : sbox_fwd = 8'h2c; 194: sbox_fwd = 8'h25;
        67 : sbox_fwd = 8'h1a; 195: sbox_fwd = 8'h2e;
        68 : sbox_fwd = 8'h1b; 196: sbox_fwd = 8'h1c;
        69 : sbox_fwd = 8'h6e; 197: sbox_fwd = 8'ha6;
        70 : sbox_fwd = 8'h5a; 198: sbox_fwd = 8'hb4;
        71 : sbox_fwd = 8'ha0; 199: sbox_fwd = 8'hc6;
        72 : sbox_fwd = 8'h52; 200: sbox_fwd = 8'he8;
        73 : sbox_fwd = 8'h3b; 201: sbox_fwd = 8'hdd;
        74 : sbox_fwd = 8'hd6; 202: sbox_fwd = 8'h74;
        75 : sbox_fwd = 8'hb3; 203: sbox_fwd = 8'h1f;
        76 : sbox_fwd = 8'h29; 204: sbox_fwd = 8'h4b;
        77 : sbox_fwd = 8'he3; 205: sbox_fwd = 8'hbd;
        78 : sbox_fwd = 8'h2f; 206: sbox_fwd = 8'h8b;
        79 : sbox_fwd = 8'h84; 207: sbox_fwd = 8'h8a;
        80 : sbox_fwd = 8'h53; 208: sbox_fwd = 8'h70;
        81 : sbox_fwd = 8'hd1; 209: sbox_fwd = 8'h3e;
        82 : sbox_fwd = 8'h00; 210: sbox_fwd = 8'hb5;
        83 : sbox_fwd = 8'hed; 211: sbox_fwd = 8'h66;
        84 : sbox_fwd = 8'h20; 212: sbox_fwd = 8'h48;
        85 : sbox_fwd = 8'hfc; 213: sbox_fwd = 8'h03;
        86 : sbox_fwd = 8'hb1; 214: sbox_fwd = 8'hf6;
        87 : sbox_fwd = 8'h5b; 215: sbox_fwd = 8'h0e;
        88 : sbox_fwd = 8'h6a; 216: sbox_fwd = 8'h61;
        89 : sbox_fwd = 8'hcb; 217: sbox_fwd = 8'h35;
        90 : sbox_fwd = 8'hbe; 218: sbox_fwd = 8'h57;
        91 : sbox_fwd = 8'h39; 219: sbox_fwd = 8'hb9;
        92 : sbox_fwd = 8'h4a; 220: sbox_fwd = 8'h86;
        93 : sbox_fwd = 8'h4c; 221: sbox_fwd = 8'hc1;
        94 : sbox_fwd = 8'h58; 222: sbox_fwd = 8'h1d;
        95 : sbox_fwd = 8'hcf; 223: sbox_fwd = 8'h9e;
        96 : sbox_fwd = 8'hd0; 224: sbox_fwd = 8'he1;
        97 : sbox_fwd = 8'hef; 225: sbox_fwd = 8'hf8;
        98 : sbox_fwd = 8'haa; 226: sbox_fwd = 8'h98;
        99 : sbox_fwd = 8'hfb; 227: sbox_fwd = 8'h11;
        100: sbox_fwd = 8'h43; 228: sbox_fwd = 8'h69;
        101: sbox_fwd = 8'h4d; 229: sbox_fwd = 8'hd9;
        102: sbox_fwd = 8'h33; 230: sbox_fwd = 8'h8e;
        103: sbox_fwd = 8'h85; 231: sbox_fwd = 8'h94;
        104: sbox_fwd = 8'h45; 232: sbox_fwd = 8'h9b;
        105: sbox_fwd = 8'hf9; 233: sbox_fwd = 8'h1e;
        106: sbox_fwd = 8'h02; 234: sbox_fwd = 8'h87;
        107: sbox_fwd = 8'h7f; 235: sbox_fwd = 8'he9;
        108: sbox_fwd = 8'h50; 236: sbox_fwd = 8'hce;
        109: sbox_fwd = 8'h3c; 237: sbox_fwd = 8'h55;
        110: sbox_fwd = 8'h9f; 238: sbox_fwd = 8'h28;
        111: sbox_fwd = 8'ha8; 239: sbox_fwd = 8'hdf;
        112: sbox_fwd = 8'h51; 240: sbox_fwd = 8'h8c;
        113: sbox_fwd = 8'ha3; 241: sbox_fwd = 8'ha1;
        114: sbox_fwd = 8'h40; 242: sbox_fwd = 8'h89;
        115: sbox_fwd = 8'h8f; 243: sbox_fwd = 8'h0d;
        116: sbox_fwd = 8'h92; 244: sbox_fwd = 8'hbf;
        117: sbox_fwd = 8'h9d; 245: sbox_fwd = 8'he6;
        118: sbox_fwd = 8'h38; 246: sbox_fwd = 8'h42;
        119: sbox_fwd = 8'hf5; 247: sbox_fwd = 8'h68;
        120: sbox_fwd = 8'hbc; 248: sbox_fwd = 8'h41;
        121: sbox_fwd = 8'hb6; 249: sbox_fwd = 8'h99;
        122: sbox_fwd = 8'hda; 250: sbox_fwd = 8'h2d;
        123: sbox_fwd = 8'h21; 251: sbox_fwd = 8'h0f;
        124: sbox_fwd = 8'h10; 252: sbox_fwd = 8'hb0;
        125: sbox_fwd = 8'hff; 253: sbox_fwd = 8'h54;
        126: sbox_fwd = 8'hf3; 254: sbox_fwd = 8'hbb;
        127: sbox_fwd = 8'hd2; 255: sbox_fwd = 8'h16;
    endcase
endfunction

//
// AES Inverse SBOX function
//
function [7:0] sbox_inv;
    input [7:0] in;

    case(in)
        0  : sbox_inv = 8'h52; 128: sbox_inv = 8'h3a;
        1  : sbox_inv = 8'h09; 129: sbox_inv = 8'h91;
        2  : sbox_inv = 8'h6a; 130: sbox_inv = 8'h11;
        3  : sbox_inv = 8'hd5; 131: sbox_inv = 8'h41;
        4  : sbox_inv = 8'h30; 132: sbox_inv = 8'h4f;
        5  : sbox_inv = 8'h36; 133: sbox_inv = 8'h67;
        6  : sbox_inv = 8'ha5; 134: sbox_inv = 8'hdc;
        7  : sbox_inv = 8'h38; 135: sbox_inv = 8'hea;
        8  : sbox_inv = 8'hbf; 136: sbox_inv = 8'h97;
        9  : sbox_inv = 8'h40; 137: sbox_inv = 8'hf2;
        10 : sbox_inv = 8'ha3; 138: sbox_inv = 8'hcf;
        11 : sbox_inv = 8'h9e; 139: sbox_inv = 8'hce;
        12 : sbox_inv = 8'h81; 140: sbox_inv = 8'hf0;
        13 : sbox_inv = 8'hf3; 141: sbox_inv = 8'hb4;
        14 : sbox_inv = 8'hd7; 142: sbox_inv = 8'he6;
        15 : sbox_inv = 8'hfb; 143: sbox_inv = 8'h73;
        16 : sbox_inv = 8'h7c; 144: sbox_inv = 8'h96;
        17 : sbox_inv = 8'he3; 145: sbox_inv = 8'hac;
        18 : sbox_inv = 8'h39; 146: sbox_inv = 8'h74;
        19 : sbox_inv = 8'h82; 147: sbox_inv = 8'h22;
        20 : sbox_inv = 8'h9b; 148: sbox_inv = 8'he7;
        21 : sbox_inv = 8'h2f; 149: sbox_inv = 8'had;
        22 : sbox_inv = 8'hff; 150: sbox_inv = 8'h35;
        23 : sbox_inv = 8'h87; 151: sbox_inv = 8'h85;
        24 : sbox_inv = 8'h34; 152: sbox_inv = 8'he2;
        25 : sbox_inv = 8'h8e; 153: sbox_inv = 8'hf9;
        26 : sbox_inv = 8'h43; 154: sbox_inv = 8'h37;
        27 : sbox_inv = 8'h44; 155: sbox_inv = 8'he8;
        28 : sbox_inv = 8'hc4; 156: sbox_inv = 8'h1c;
        29 : sbox_inv = 8'hde; 157: sbox_inv = 8'h75;
        30 : sbox_inv = 8'he9; 158: sbox_inv = 8'hdf;
        31 : sbox_inv = 8'hcb; 159: sbox_inv = 8'h6e;
        32 : sbox_inv = 8'h54; 160: sbox_inv = 8'h47;
        33 : sbox_inv = 8'h7b; 161: sbox_inv = 8'hf1;
        34 : sbox_inv = 8'h94; 162: sbox_inv = 8'h1a;
        35 : sbox_inv = 8'h32; 163: sbox_inv = 8'h71;
        36 : sbox_inv = 8'ha6; 164: sbox_inv = 8'h1d;
        37 : sbox_inv = 8'hc2; 165: sbox_inv = 8'h29;
        38 : sbox_inv = 8'h23; 166: sbox_inv = 8'hc5;
        39 : sbox_inv = 8'h3d; 167: sbox_inv = 8'h89;
        40 : sbox_inv = 8'hee; 168: sbox_inv = 8'h6f;
        41 : sbox_inv = 8'h4c; 169: sbox_inv = 8'hb7;
        42 : sbox_inv = 8'h95; 170: sbox_inv = 8'h62;
        43 : sbox_inv = 8'h0b; 171: sbox_inv = 8'h0e;
        44 : sbox_inv = 8'h42; 172: sbox_inv = 8'haa;
        45 : sbox_inv = 8'hfa; 173: sbox_inv = 8'h18;
        46 : sbox_inv = 8'hc3; 174: sbox_inv = 8'hbe;
        47 : sbox_inv = 8'h4e; 175: sbox_inv = 8'h1b;
        48 : sbox_inv = 8'h08; 176: sbox_inv = 8'hfc;
        49 : sbox_inv = 8'h2e; 177: sbox_inv = 8'h56;
        50 : sbox_inv = 8'ha1; 178: sbox_inv = 8'h3e;
        51 : sbox_inv = 8'h66; 179: sbox_inv = 8'h4b;
        52 : sbox_inv = 8'h28; 180: sbox_inv = 8'hc6;
        53 : sbox_inv = 8'hd9; 181: sbox_inv = 8'hd2;
        54 : sbox_inv = 8'h24; 182: sbox_inv = 8'h79;
        55 : sbox_inv = 8'hb2; 183: sbox_inv = 8'h20;
        56 : sbox_inv = 8'h76; 184: sbox_inv = 8'h9a;
        57 : sbox_inv = 8'h5b; 185: sbox_inv = 8'hdb;
        58 : sbox_inv = 8'ha2; 186: sbox_inv = 8'hc0;
        59 : sbox_inv = 8'h49; 187: sbox_inv = 8'hfe;
        60 : sbox_inv = 8'h6d; 188: sbox_inv = 8'h78;
        61 : sbox_inv = 8'h8b; 189: sbox_inv = 8'hcd;
        62 : sbox_inv = 8'hd1; 190: sbox_inv = 8'h5a;
        63 : sbox_inv = 8'h25; 191: sbox_inv = 8'hf4;
        64 : sbox_inv = 8'h72; 192: sbox_inv = 8'h1f;
        65 : sbox_inv = 8'hf8; 193: sbox_inv = 8'hdd;
        66 : sbox_inv = 8'hf6; 194: sbox_inv = 8'ha8;
        67 : sbox_inv = 8'h64; 195: sbox_inv = 8'h33;
        68 : sbox_inv = 8'h86; 196: sbox_inv = 8'h88;
        69 : sbox_inv = 8'h68; 197: sbox_inv = 8'h07;
        70 : sbox_inv = 8'h98; 198: sbox_inv = 8'hc7;
        71 : sbox_inv = 8'h16; 199: sbox_inv = 8'h31;
        72 : sbox_inv = 8'hd4; 200: sbox_inv = 8'hb1;
        73 : sbox_inv = 8'ha4; 201: sbox_inv = 8'h12;
        74 : sbox_inv = 8'h5c; 202: sbox_inv = 8'h10;
        75 : sbox_inv = 8'hcc; 203: sbox_inv = 8'h59;
        76 : sbox_inv = 8'h5d; 204: sbox_inv = 8'h27;
        77 : sbox_inv = 8'h65; 205: sbox_inv = 8'h80;
        78 : sbox_inv = 8'hb6; 206: sbox_inv = 8'hec;
        79 : sbox_inv = 8'h92; 207: sbox_inv = 8'h5f;
        80 : sbox_inv = 8'h6c; 208: sbox_inv = 8'h60;
        81 : sbox_inv = 8'h70; 209: sbox_inv = 8'h51;
        82 : sbox_inv = 8'h48; 210: sbox_inv = 8'h7f;
        83 : sbox_inv = 8'h50; 211: sbox_inv = 8'ha9;
        84 : sbox_inv = 8'hfd; 212: sbox_inv = 8'h19;
        85 : sbox_inv = 8'hed; 213: sbox_inv = 8'hb5;
        86 : sbox_inv = 8'hb9; 214: sbox_inv = 8'h4a;
        87 : sbox_inv = 8'hda; 215: sbox_inv = 8'h0d;
        88 : sbox_inv = 8'h5e; 216: sbox_inv = 8'h2d;
        89 : sbox_inv = 8'h15; 217: sbox_inv = 8'he5;
        90 : sbox_inv = 8'h46; 218: sbox_inv = 8'h7a;
        91 : sbox_inv = 8'h57; 219: sbox_inv = 8'h9f;
        92 : sbox_inv = 8'ha7; 220: sbox_inv = 8'h93;
        93 : sbox_inv = 8'h8d; 221: sbox_inv = 8'hc9;
        94 : sbox_inv = 8'h9d; 222: sbox_inv = 8'h9c;
        95 : sbox_inv = 8'h84; 223: sbox_inv = 8'hef;
        96 : sbox_inv = 8'h90; 224: sbox_inv = 8'ha0;
        97 : sbox_inv = 8'hd8; 225: sbox_inv = 8'he0;
        98 : sbox_inv = 8'hab; 226: sbox_inv = 8'h3b;
        99 : sbox_inv = 8'h00; 227: sbox_inv = 8'h4d;
        100: sbox_inv = 8'h8c; 228: sbox_inv = 8'hae;
        101: sbox_inv = 8'hbc; 229: sbox_inv = 8'h2a;
        102: sbox_inv = 8'hd3; 230: sbox_inv = 8'hf5;
        103: sbox_inv = 8'h0a; 231: sbox_inv = 8'hb0;
        104: sbox_inv = 8'hf7; 232: sbox_inv = 8'hc8;
        105: sbox_inv = 8'he4; 233: sbox_inv = 8'heb;
        106: sbox_inv = 8'h58; 234: sbox_inv = 8'hbb;
        107: sbox_inv = 8'h05; 235: sbox_inv = 8'h3c;
        108: sbox_inv = 8'hb8; 236: sbox_inv = 8'h83;
        109: sbox_inv = 8'hb3; 237: sbox_inv = 8'h53;
        110: sbox_inv = 8'h45; 238: sbox_inv = 8'h99;
        111: sbox_inv = 8'h06; 239: sbox_inv = 8'h61;
        112: sbox_inv = 8'hd0; 240: sbox_inv = 8'h17;
        113: sbox_inv = 8'h2c; 241: sbox_inv = 8'h2b;
        114: sbox_inv = 8'h1e; 242: sbox_inv = 8'h04;
        115: sbox_inv = 8'h8f; 243: sbox_inv = 8'h7e;
        116: sbox_inv = 8'hca; 244: sbox_inv = 8'hba;
        117: sbox_inv = 8'h3f; 245: sbox_inv = 8'h77;
        118: sbox_inv = 8'h0f; 246: sbox_inv = 8'hd6;
        119: sbox_inv = 8'h02; 247: sbox_inv = 8'h26;
        120: sbox_inv = 8'hc1; 248: sbox_inv = 8'he1;
        121: sbox_inv = 8'haf; 249: sbox_inv = 8'h69;
        122: sbox_inv = 8'hbd; 250: sbox_inv = 8'h14;
        123: sbox_inv = 8'h03; 251: sbox_inv = 8'h63;
        124: sbox_inv = 8'h01; 252: sbox_inv = 8'h55;
        125: sbox_inv = 8'h13; 253: sbox_inv = 8'h21;
        126: sbox_inv = 8'h8a; 254: sbox_inv = 8'h0c;
        127: sbox_inv = 8'h6b; 255: sbox_inv = 8'h7d;
    endcase
endfunction
