//
// SCARV Project
// 
// University of Bristol
// 
// RISC-V Cryptographic Instruction Set Extension
// 
// Reference Implementation
// 
// 

//
// module: tb_formal
//
//  Top level testbench for the formal verification flow.
//
module tb_formal ();




endmodule

